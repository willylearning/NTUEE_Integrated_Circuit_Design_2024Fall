* File: adder.pex.sp
* Created: Fri Nov  8 13:28:07 2024
* Program "Calibre xRC"
* Version "v2022.3_33.19"
* 
.include "adder.pex.sp.pex"
.subckt adder  S1 S2 S3 COUT S4 A1 VDD GND B1 CIN C1 A2 B2 C2 A3 C3 A4 B4
* 
* B4	B4
* A4	A4
* C3	C3
* A3	A3
* C2	C2
* B2	B2
* A2	A2
* C1	C1
* CIN	CIN
* B1	B1
* GND	GND
* VDD	VDD
* A1	A1
* S4	S4
* COUT	COUT
* S3	S3
* S2	S2
* S1	S1
M5 N_D3_M5_d N_A1_M5_g N_GND_M5_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06 AD=8.2e-13
+ AS=8e-13 PD=2.64e-06 PS=2.6e-06
M6 N_D3_M6_d N_B1_M6_g N_GND_M6_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06 AD=8.2e-13
+ AS=8e-13 PD=2.64e-06 PS=2.6e-06
M4 N_D2_M4_d N_CIN_M4_g N_D3_M4_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06 AD=8.2e-13
+ AS=8e-13 PD=2.64e-06 PS=2.6e-06
M10 N_D5_M10_d N_A1_M10_g N_GND_M10_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M9 N_D2_M9_d N_B1_M9_g N_D5_M9_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06 AD=8.2e-13
+ AS=8e-13 PD=2.64e-06 PS=2.6e-06
M26 N_C1_M26_d N_D2_M26_g N_GND_M26_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M16 N_D8_M16_d N_A1_M16_g N_GND_M16_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M17 N_D8_M17_d N_B1_M17_g N_GND_M17_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M18 N_D8_M18_d N_CIN_M18_g N_GND_M18_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M15 N_D7_M15_d N_D2_M15_g N_D8_M15_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M24 N_D12_M24_d N_A1_M24_g N_GND_M24_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M23 N_D11_M23_d N_B1_M23_g N_D12_M23_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M22 N_D7_M22_d N_CIN_M22_g N_D11_M22_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M28 N_S1_M28_d N_D7_M28_g N_GND_M28_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M33 N_E3_M33_d N_A2_M33_g N_GND_M33_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M34 N_E3_M34_d N_B2_M34_g N_GND_M34_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M32 N_E2_M32_d N_C1_M32_g N_E3_M32_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M38 N_E5_M38_d N_A2_M38_g N_GND_M38_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M37 N_E2_M37_d N_B2_M37_g N_E5_M37_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M54 N_C2_M54_d N_E2_M54_g N_GND_M54_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M44 N_E8_M44_d N_A2_M44_g N_GND_M44_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M45 N_E8_M45_d N_B2_M45_g N_GND_M45_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M46 N_E8_M46_d N_C1_M46_g N_GND_M46_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M43 N_E7_M43_d N_E2_M43_g N_E8_M43_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M52 N_E12_M52_d N_A2_M52_g N_GND_M52_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M51 N_E11_M51_d N_B2_M51_g N_E12_M51_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M50 N_E7_M50_d N_C1_M50_g N_E11_M50_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M56 N_S2_M56_d N_E7_M56_g N_GND_M56_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M61 N_F3_M61_d N_A3_M61_g N_GND_M61_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M62 N_F3_M62_d N_B3_M62_g N_GND_M62_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M60 N_F2_M60_d N_C2_M60_g N_F3_M60_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M66 N_F5_M66_d N_A3_M66_g N_GND_M66_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M65 N_F2_M65_d N_B3_M65_g N_F5_M65_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M82 N_C3_M82_d N_F2_M82_g N_GND_M82_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M72 N_F8_M72_d N_A3_M72_g N_GND_M72_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M73 N_F8_M73_d N_B3_M73_g N_GND_M73_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M74 N_F8_M74_d N_C2_M74_g N_GND_M74_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M71 N_F7_M71_d N_F2_M71_g N_F8_M71_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M80 N_F12_M80_d N_A3_M80_g N_GND_M80_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M79 N_F11_M79_d N_B3_M79_g N_F12_M79_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M78 N_F7_M78_d N_C2_M78_g N_F11_M78_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M84 N_S3_M84_d N_F7_M84_g N_GND_M84_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M89 N_G3_M89_d N_A4_M89_g N_GND_M89_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M90 N_G3_M90_d N_B4_M90_g N_GND_M90_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M88 N_G2_M88_d N_C3_M88_g N_G3_M88_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M94 N_G5_M94_d N_A4_M94_g N_GND_M94_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M93 N_G2_M93_d N_B4_M93_g N_G5_M93_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M110 N_COUT_M110_d N_G2_M110_g N_GND_M110_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M100 N_G8_M100_d N_A4_M100_g N_GND_M100_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M101 N_G8_M101_d N_B4_M101_g N_GND_M101_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M102 N_G8_M102_d N_C3_M102_g N_GND_M102_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M99 N_G7_M99_d N_G2_M99_g N_G8_M99_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M108 N_G12_M108_d N_A4_M108_g N_GND_M108_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M107 N_G11_M107_d N_B4_M107_g N_G12_M107_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M106 N_G7_M106_d N_C3_M106_g N_G11_M106_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M112 N_S4_M112_d N_G7_M112_g N_GND_M112_s N_GND_M5_b N_18 L=1.8e-07 W=1e-06
+ AD=8.2e-13 AS=8e-13 PD=2.64e-06 PS=2.6e-06
M1 N_D1_M1_d N_A1_M1_g N_VDD_M1_s N_VDD_M1_b P_18 L=1.8e-07 W=2e-06 AD=1.64e-12
+ AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M2 N_D1_M2_d N_B1_M2_g N_VDD_M2_s N_VDD_M2_b P_18 L=1.8e-07 W=2e-06 AD=1.64e-12
+ AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M3 N_D2_M3_d N_CIN_M3_g N_D1_M3_s N_VDD_M3_b P_18 L=1.8e-07 W=2e-06 AD=1.64e-12
+ AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M7 N_D4_M7_d N_A1_M7_g N_VDD_M7_s N_VDD_M7_b P_18 L=1.8e-07 W=2e-06 AD=1.64e-12
+ AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M8 N_D2_M8_d N_B1_M8_g N_D4_M8_s N_VDD_M8_b P_18 L=1.8e-07 W=2e-06 AD=1.64e-12
+ AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M25 N_C1_M25_d N_D2_M25_g N_VDD_M25_s N_VDD_M25_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M13 N_D6_M13_d N_CIN_M13_g N_VDD_M13_s N_VDD_M13_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M12 N_D6_M12_d N_B1_M12_g N_VDD_M12_s N_VDD_M12_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M11 N_D6_M11_d N_A1_M11_g N_VDD_M11_s N_VDD_M11_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M14 N_D7_M14_d N_D2_M14_g N_D6_M14_s N_VDD_M14_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M19 N_D9_M19_d N_A1_M19_g N_VDD_M19_s N_VDD_M19_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M20 N_D10_M20_d N_B1_M20_g N_D9_M20_s N_VDD_M20_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M21 N_D7_M21_d N_CIN_M21_g N_D10_M21_s N_VDD_M21_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M27 N_S1_M27_d N_D7_M27_g N_VDD_M27_s N_VDD_M27_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M29 N_E1_M29_d N_A2_M29_g N_VDD_M29_s N_VDD_M29_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M30 N_E1_M30_d N_B2_M30_g N_VDD_M30_s N_VDD_M30_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M31 N_E2_M31_d N_C1_M31_g N_E1_M31_s N_VDD_M31_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M35 N_E4_M35_d N_A2_M35_g N_VDD_M35_s N_VDD_M35_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M36 N_E2_M36_d N_B2_M36_g N_E4_M36_s N_VDD_M36_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M53 N_C2_M53_d N_E2_M53_g N_VDD_M53_s N_VDD_M53_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M41 N_E6_M41_d N_C1_M41_g N_VDD_M41_s N_VDD_M41_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M40 N_E6_M40_d N_B2_M40_g N_VDD_M40_s N_VDD_M40_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M39 N_E6_M39_d N_A2_M39_g N_VDD_M39_s N_VDD_M39_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M42 N_E7_M42_d N_E2_M42_g N_E6_M42_s N_VDD_M42_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M47 N_E9_M47_d N_A2_M47_g N_VDD_M47_s N_VDD_M47_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M48 N_E10_M48_d N_B2_M48_g N_E9_M48_s N_VDD_M48_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M49 N_E7_M49_d N_C1_M49_g N_E10_M49_s N_VDD_M49_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M55 N_S2_M55_d N_E7_M55_g N_VDD_M55_s N_VDD_M55_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M57 N_F1_M57_d N_A3_M57_g N_VDD_M57_s N_VDD_M57_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M58 N_F1_M58_d N_B3_M58_g N_VDD_M58_s N_VDD_M58_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M59 N_F2_M59_d N_C2_M59_g N_F1_M59_s N_VDD_M59_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M63 N_F4_M63_d N_A3_M63_g N_VDD_M63_s N_VDD_M63_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M64 N_F2_M64_d N_B3_M64_g N_F4_M64_s N_VDD_M64_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M81 N_C3_M81_d N_F2_M81_g N_VDD_M81_s N_VDD_M81_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M69 N_F6_M69_d N_C2_M69_g N_VDD_M69_s N_VDD_M69_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M68 N_F6_M68_d N_B3_M68_g N_VDD_M68_s N_VDD_M68_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M67 N_F6_M67_d N_A3_M67_g N_VDD_M67_s N_VDD_M67_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M70 N_F7_M70_d N_F2_M70_g N_F6_M70_s N_VDD_M70_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M75 N_F9_M75_d N_A3_M75_g N_VDD_M75_s N_VDD_M75_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M76 N_F10_M76_d N_B3_M76_g N_F9_M76_s N_VDD_M76_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M77 N_F7_M77_d N_C2_M77_g N_F10_M77_s N_VDD_M77_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M83 N_S3_M83_d N_F7_M83_g N_VDD_M83_s N_VDD_M83_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M85 N_G1_M85_d N_A4_M85_g N_VDD_M85_s N_VDD_M85_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M86 N_G1_M86_d N_B4_M86_g N_VDD_M86_s N_VDD_M86_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M87 N_G2_M87_d N_C3_M87_g N_G1_M87_s N_VDD_M87_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M91 N_G4_M91_d N_A4_M91_g N_VDD_M91_s N_VDD_M91_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M92 N_G2_M92_d N_B4_M92_g N_G4_M92_s N_VDD_M92_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M109 N_COUT_M109_d N_G2_M109_g N_VDD_M109_s N_VDD_M109_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M97 N_G6_M97_d N_C3_M97_g N_VDD_M97_s N_VDD_M97_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M96 N_G6_M96_d N_B4_M96_g N_VDD_M96_s N_VDD_M96_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M95 N_G6_M95_d N_A4_M95_g N_VDD_M95_s N_VDD_M95_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M98 N_G7_M98_d N_G2_M98_g N_G6_M98_s N_VDD_M98_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M103 N_G9_M103_d N_A4_M103_g N_VDD_M103_s N_VDD_M103_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M104 N_G10_M104_d N_B4_M104_g N_G9_M104_s N_VDD_M104_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M105 N_G7_M105_d N_C3_M105_g N_G10_M105_s N_VDD_M105_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
M111 N_S4_M111_d N_G7_M111_g N_VDD_M111_s N_VDD_M111_b P_18 L=1.8e-07 W=2e-06
+ AD=1.64e-12 AS=1.6e-12 PD=3.64e-06 PS=3.6e-06
*
.include "adder.pex.sp.ADDER.pxi"
*
.ends
*
*
